module MXU (
    input [143:0] A,
    input [143:0] B,
    output [143:0] mxu_out
);

    assign mxu_out = {
        {A[111:96] * B[47:32] + A[127:112] * B[95:80] + A[143:128] * B[143:128]},
        {A[111:96] * B[31:16] + A[127:112] * B[79:64] + A[143:128] * B[127:112]},
        {A[111:96] * B[15:0] + A[127:112] * B[63:48] + A[143:128] * B[111:96]},
        {A[63:48] * B[47:32] + A[79:64] * B[95:80] + A[95:80] * B[143:128]},
        {A[63:48] * B[31:16] + A[79:64] * B[79:64] + A[95:80] * B[127:112]},
        {A[63:48] * B[15:0] + A[79:64] * B[63:48] + A[95:80] * B[111:96]},
        {A[15:0] * B[47:32] + A[31:16] * B[95:80] + A[47:32] * B[143:128]},
        {A[15:0] * B[31:16] + A[31:16] * B[79:64] + A[47:32] * B[127:112]},
        {A[15:0] * B[15:0] + A[31:16] * B[63:48] + A[47:32] * B[111:96]}
    };

endmodule